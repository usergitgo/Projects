`timescale 1ns / 1ps

module Cartoon_Filter #(  // Gaussian blur -> posterize -> Sobel edge overlay
    parameter int IMG_WIDTH    = 320,
    parameter int IMG_HEIGHT   = 240,
    // Posterization level (keep MSBs)
    parameter int KEEP_RB_MSBS = 2,    // 1..5 (R/B 5bit)
    parameter int KEEP_G_MSBS  = 2,    // 1..6 (G  6bit)
    // Edge threshold (|Gx|+|Gy|)
    parameter int EDGE_THR     = 50
) (
    input logic        clk,
    input logic        reset,
    // camera write stream
    input logic        we_in,
    input logic [16:0] wAddr_in,
    input logic [15:0] wData_in,

    // to frame buffer
    output logic        we_out,
    output logic [16:0] wAddr_out,
    output logic [15:0] wData_out
);

    // ---------------------------------------------------------
    // 1) Coordinate counters
    // ---------------------------------------------------------
    logic [$clog2(IMG_WIDTH )-1:0] col_cnt;
    logic [$clog2(IMG_HEIGHT)-1:0] row_cnt;
    wire frame_start = (we_in && (wAddr_in == 17'd0));

    always_ff @(posedge clk) begin
        if (reset) begin
            col_cnt <= '0;
            row_cnt <= '0;
        end else if (we_in) begin
            if (frame_start) begin
                col_cnt <= '0;
                row_cnt <= '0;
            end else if (col_cnt == IMG_WIDTH - 1) begin
                col_cnt <= '0;
                row_cnt <= (row_cnt == IMG_HEIGHT - 1) ? '0 : (row_cnt + 1'b1);
            end else begin
                col_cnt <= col_cnt + 1'b1;
            end
        end
    end

    // ---------------------------------------------------------
    // 2) RGB565 split
    // ---------------------------------------------------------
    logic [4:0] in_r5;
    logic [5:0] in_g6;
    logic [4:0] in_b5;
    always_comb begin
        in_r5 = wData_in[15:11];
        in_g6 = wData_in[10:5];
        in_b5 = wData_in[4:0];
    end

    // ---------------------------------------------------------
    // 3) Line buffers + 3x3 window
    // ---------------------------------------------------------
    logic [4:0] line1_r[0:IMG_WIDTH-1], line2_r[0:IMG_WIDTH-1];
    logic [5:0] line1_g[0:IMG_WIDTH-1], line2_g[0:IMG_WIDTH-1];
    logic [4:0] line1_b[0:IMG_WIDTH-1], line2_b[0:IMG_WIDTH-1];

    logic [4:0] r00, r01, r02, r10, r11, r12, r20, r21, r22;
    logic [5:0] g00, g01, g02, g10, g11, g12, g20, g21, g22;
    logic [4:0] b00, b01, b02, b10, b11, b12, b20, b21, b22;

    logic [15:0] raw_pixel_d1, raw_pixel_d2;
    logic [16:0] addr_d1, addr_d2, addr_d3;
    logic we_d1, we_d2, we_d3;

    wire  at_border_now = (col_cnt==0) || (row_cnt==0)
                       || (col_cnt==IMG_WIDTH-1) || (row_cnt==IMG_HEIGHT-1);
    logic at_border_d1, at_border_d2;

    always_ff @(posedge clk) begin
        if (reset) begin
            {r00, r01, r02, r10, r11, r12, r20, r21, r22} <= '{default: '0};
            {g00, g01, g02, g10, g11, g12, g20, g21, g22} <= '{default: '0};
            {b00, b01, b02, b10, b11, b12, b20, b21, b22} <= '{default: '0};
            raw_pixel_d1 <= '0;
            raw_pixel_d2 <= '0;
            addr_d1 <= '0;
            addr_d2 <= '0;
            addr_d3 <= '0;
            we_d1 <= 1'b0;
            we_d2 <= 1'b0;
            we_d3 <= 1'b0;
            at_border_d1 <= 1'b0;
            at_border_d2 <= 1'b0;
        end else begin
            raw_pixel_d1 <= wData_in;
            raw_pixel_d2 <= raw_pixel_d1;
            addr_d1 <= wAddr_in;
            addr_d2 <= addr_d1;
            addr_d3 <= addr_d2;
            we_d1 <= we_in;
            we_d2 <= we_d1;
            we_d3 <= we_d2;
            at_border_d1 <= at_border_now;
            at_border_d2 <= at_border_d1;

            if (we_in) begin
                r00 <= r01;
                r01 <= r02;
                r02 <= line2_r[col_cnt];
                r10 <= r11;
                r11 <= r12;
                r12 <= line1_r[col_cnt];
                r20 <= r21;
                r21 <= r22;
                r22 <= in_r5;

                g00 <= g01;
                g01 <= g02;
                g02 <= line2_g[col_cnt];
                g10 <= g11;
                g11 <= g12;
                g12 <= line1_g[col_cnt];
                g20 <= g21;
                g21 <= g22;
                g22 <= in_g6;

                b00 <= b01;
                b01 <= b02;
                b02 <= line2_b[col_cnt];
                b10 <= b11;
                b11 <= b12;
                b12 <= line1_b[col_cnt];
                b20 <= b21;
                b21 <= b22;
                b22 <= in_b5;

                line2_r[col_cnt] <= line1_r[col_cnt];
                line1_r[col_cnt] <= in_r5;
                line2_g[col_cnt] <= line1_g[col_cnt];
                line1_g[col_cnt] <= in_g6;
                line2_b[col_cnt] <= line1_b[col_cnt];
                line1_b[col_cnt] <= in_b5;
            end
        end
    end

    // ---------------------------------------------------------
    // 4) 3x3 Gaussian blur (1 2 1; 2 4 2; 1 2 1)/16
    // ---------------------------------------------------------
    logic [11:0] sum_r, sum_g, sum_b;
    logic [4:0] blur_r5;
    logic [5:0] blur_g6;
    logic [4:0] blur_b5;

    always_ff @(posedge clk) begin
        if (reset) begin
            sum_r   <= '0;
            sum_g   <= '0;
            sum_b   <= '0;
            blur_r5 <= '0;
            blur_g6 <= '0;
            blur_b5 <= '0;
        end else begin
            sum_r <= (r00 + (r01<<1) + r02)
                   + ((r10<<1) + (r11<<2) + (r12<<1))
                   + (r20 + (r21<<1) + r22);
            sum_g <= (g00 + (g01<<1) + g02)
                   + ((g10<<1) + (g11<<2) + (g12<<1))
                   + (g20 + (g21<<1) + g22);
            sum_b <= (b00 + (b01<<1) + b02)
                   + ((b10<<1) + (b11<<2) + (b12<<1))
                   + (b20 + (b21<<1) + b22);

            blur_r5 <= (sum_r[11:4] > 12'd31) ? 5'd31 : sum_r[8:4];
            blur_g6 <= (sum_g[11:4] > 12'd63) ? 6'd63 : sum_g[9:4];
            blur_b5 <= (sum_b[11:4] > 12'd31) ? 5'd31 : sum_b[8:4];
        end
    end

    // ---------------------------------------------------------
    // 5) Posterization (keep MSBs, zero LSBs) — generate-if로 분기
    // ---------------------------------------------------------
    wire [4:0] post_r5_w;
    wire [5:0] post_g6_w;
    wire [4:0] post_b5_w;

    generate
        if (KEEP_RB_MSBS >= 5) begin
            assign post_r5_w = blur_r5;
            assign post_b5_w = blur_b5;
        end else if (KEEP_RB_MSBS == 4) begin
            assign post_r5_w = {blur_r5[4:1], 1'b0};
            assign post_b5_w = {blur_b5[4:1], 1'b0};
        end else if (KEEP_RB_MSBS == 3) begin
            assign post_r5_w = {blur_r5[4:2], 2'b00};
            assign post_b5_w = {blur_b5[4:2], 2'b00};
        end else if (KEEP_RB_MSBS == 2) begin
            assign post_r5_w = {blur_r5[4:3], 3'b000};
            assign post_b5_w = {blur_b5[4:3], 3'b000};
        end else begin  // KEEP_RB_MSBS == 1 (or less)
            assign post_r5_w = {blur_r5[4], 4'b0000};
            assign post_b5_w = {blur_b5[4], 4'b0000};
        end
    endgenerate

    generate
        if (KEEP_G_MSBS >= 6) begin
            assign post_g6_w = blur_g6;
        end else if (KEEP_G_MSBS == 5) begin
            assign post_g6_w = {blur_g6[5:1], 1'b0};
        end else if (KEEP_G_MSBS == 4) begin
            assign post_g6_w = {blur_g6[5:2], 2'b00};
        end else if (KEEP_G_MSBS == 3) begin
            assign post_g6_w = {blur_g6[5:3], 3'b000};
        end else if (KEEP_G_MSBS == 2) begin
            assign post_g6_w = {blur_g6[5:4], 4'b0000};
        end else begin  // KEEP_G_MSBS == 1 (or less)
            assign post_g6_w = {blur_g6[5], 5'b00000};
        end
    endgenerate

    logic [4:0] post_r5;
    logic [5:0] post_g6;
    logic [4:0] post_b5;
    always_ff @(posedge clk) begin
        if (reset) begin
            post_r5 <= '0;
            post_g6 <= '0;
            post_b5 <= '0;
        end else begin
            post_r5 <= post_r5_w;
            post_g6 <= post_g6_w;
            post_b5 <= post_b5_w;
        end
    end

    // ---------------------------------------------------------
    // 6) Sobel edge on G (|Gx| + |Gy|)
    // ---------------------------------------------------------
    logic signed [10:0] gx, gy;
    logic [10:0] abs_gx, abs_gy;
    logic [11:0] edge_mag;

    always_ff @(posedge clk) begin
        if (reset) begin
            gx <= '0;
            gy <= '0;
            abs_gx <= '0;
            abs_gy <= '0;
            edge_mag <= '0;
        end else begin
            gx <= $signed(
                {1'b0, g02}
            ) + $signed(
                {1'b0, (g12 << 1)}
            ) + $signed(
                {1'b0, g22}
            ) - ($signed(
                {1'b0, g00}
            ) + $signed(
                {1'b0, (g10 << 1)}
            ) + $signed(
                {1'b0, g20}
            ));
            gy <= $signed(
                {1'b0, g20}
            ) + $signed(
                {1'b0, (g21 << 1)}
            ) + $signed(
                {1'b0, g22}
            ) - ($signed(
                {1'b0, g00}
            ) + $signed(
                {1'b0, (g01 << 1)}
            ) + $signed(
                {1'b0, g02}
            ));

            abs_gx <= gx[10] ? (~gx + 11'd1) : gx;
            abs_gy <= gy[10] ? (~gy + 11'd1) : gy;
            edge_mag <= abs_gx + abs_gy;
        end
    end

    // ---------------------------------------------------------
    // 7) Border passthrough / Edge overlay / Pack
    // ---------------------------------------------------------
    logic [4:0] out_r5;
    logic [5:0] out_g6;
    logic [4:0] out_b5;

    always_ff @(posedge clk) begin
        if (reset) begin
            out_r5 <= '0;
            out_g6 <= '0;
            out_b5 <= '0;
        end else if (at_border_d2) begin
            out_r5 <= raw_pixel_d2[15:11];
            out_g6 <= raw_pixel_d2[10:5];
            out_b5 <= raw_pixel_d2[4:0];
        end else begin
            if (edge_mag >= EDGE_THR) begin
                out_r5 <= 5'd0;
                out_g6 <= 6'd0;
                out_b5 <= 5'd0;  // black edge
            end else begin
                out_r5 <= post_r5;
                out_g6 <= post_g6;
                out_b5 <= post_b5;  // flat color
            end
        end
    end

    assign wData_out = {out_r5, out_g6, out_b5};

    // ---------------------------------------------------------
    // 8) Output timing
    // ---------------------------------------------------------
    always_ff @(posedge clk) begin
        if (reset) begin
            wAddr_out <= '0;
            we_out <= 1'b0;
        end else begin
            wAddr_out <= addr_d3;
            we_out    <= we_d3;
        end
    end

endmodule
